`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:24:01 04/29/2013 
// Design Name: 
// Module Name:    mode_generator 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mode_generator(
    input clk_in,
    input reset,
    output pan_pause,
    output tilt_pause,
    output pan_load,
    output tilt_load,
    output [7:0] pan_load_vec,
    output [7:0] tilt_load_vec,
    input [3:0] mode_sel
    );


endmodule
